module lab4iramHRMmod(CLK, RESET, ADDR, Q);
  input         CLK;
  input         RESET;
  input  [7:0]  ADDR;
  output [15:0] Q;

  reg    [15:0] mem[0:127]; // instruction memory with 16 bit entries

  wire   [6:0]  saddr;
  integer       i;

  assign saddr = ADDR[7:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
    if(RESET) begin

      // data goes here
      mem[0] <= 16'b1111000000000001; //   SUB R0, R0, R0
      mem[1] <= 16'b1111010010010001; //   SUB R2, R2, R2
      mem[2] <= 16'b1111111111111001; //   SUB R7, R7, R7
      mem[3] <= 16'b1111110110110001; //   SUB R6, R6, R6
      mem[4] <= 16'b0101000101111111; //   ADDI R5, R0, -1
      mem[5] <= 16'b1111101000101011; //   SRL R5, R5
      mem[6] <= 16'b0010000011111011; //   LB R3, -5(R0)
      mem[7] <= 16'b0110011011000001; //   ANDI R3, R3, 1
      mem[8] <= 16'b0010000100111011; //   LB R4, -5(R0)
      mem[9] <= 16'b0110100100000001; //   ANDI R4, R4, 1
      mem[10] <= 16'b1111100011011000; //   ADD R3, R4, R3
      mem[11] <= 16'b0110011011000001; //   ANDI R3, R3, 1
      mem[12] <= 16'b1111011100011101; //   AND R3, R3, R4
      mem[13] <= 16'b1111010011010000; //   ADD R2, R2, R3
      mem[14] <= 16'b1111100000011000; //   ADD R3, R4, R0
      mem[15] <= 16'b0101111111111111; //   ADDI R7, R7, -1
      mem[16] <= 16'b1001000111110111; //   BNE R7, R0, -9
      mem[17] <= 16'b0101110110111111; //   ADDI R6, R6, -1
      mem[18] <= 16'b1001000110110101; //   BNE R6, R0, -11
      mem[19] <= 16'b0101101101111111; //   ADDI R5, R5, -1
      mem[20] <= 16'b1001000101110011; //   BNE R5, R0, -13
      mem[21] <= 16'b0101010100100010; //   ADDI R4, R2, -30
      mem[22] <= 16'b1011100000000001; //   BLTZ R4, 1
      mem[23] <= 16'b0101000010011101; //   ADDI R2, R0, 29
      mem[24] <= 16'b1111010000010100; //   SLL R2, R2
      mem[25] <= 16'b0010010011000000; //   LB R3, 0(R2)
      mem[26] <= 16'b0100000011111110; //   SB R3, -2(R0)
      mem[27] <= 16'b0010010011000001; //   LB R3, 1(R2)
      mem[28] <= 16'b0100000011111111; //   SB R3, -1(R0)
      mem[29] <= 16'b0101111011000000; //   ADDI R3, R7, 0
      mem[30] <= 16'b1111110110110001; //   SUB R6, R6, R6
      mem[31] <= 16'b1111010000010010; //   SRA R2,R2
      mem[32] <= 16'b1001000001000001; //   BNE R1, R0, 1
      mem[33] <= 16'b0010000001111001; //   LB R1, -7(R0)
      mem[34] <= 16'b1001000101000001; //   BNE R5, R0, 1
      mem[35] <= 16'b1111010101101000; //   ADD R5, R2, R5
      mem[36] <= 16'b1000010101010011; //   BEQ R5, R2, 19
      mem[37] <= 16'b1111101010111001; //   SUB R7, R5, R2
      mem[38] <= 16'b1011111000000001; //   BLTZ R7,1
      mem[39] <= 16'b1010111000000101; //   BGEZ R7, 5
      mem[40] <= 16'b1111111001111000; //   ADD R7, R7, R1
      mem[41] <= 16'b1010111000001111; //   BGEZ R7, 15
      mem[42] <= 16'b1111111111111001; //   SUB R7, R7, R7
      mem[43] <= 16'b1000111011010000; //   BEQ R3, R7, 16
      mem[44] <= 16'b1001111011000100; //   BNE R3, R7, 4
      mem[45] <= 16'b1111111001111001; //   SUB R7, R7, R1
      mem[46] <= 16'b1011111000001100; //   BLTZ R7, 12
      mem[47] <= 16'b0101000111000001; //   ADDI R7, R0, 1
      mem[48] <= 16'b1000111011000111; //   BEQ R3, R7, 7
      mem[49] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[50] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[51] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[52] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[53] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[54] <= 16'b0101110110011001; //   ADDI R6, R6, 25
      mem[55] <= 16'b0101110110010100; //   ADDI R6, R6, 20
      mem[56] <= 16'b1011110000000011; //   BLTZ R6, 3
      mem[57] <= 16'b1111111111111001; //   SUB R7, R7, R7
      mem[58] <= 16'b1000000111000001; //   BEQ R7, R0, 1
      mem[59] <= 16'b0101000111000001; //   ADDI R7, R0, 1
      mem[60] <= 16'b0100000110111101; //   SB R6, -3(R0)
      mem[61] <= 16'b1111010000101000; //   ADD R5, R2, R0

      for(i = 62; i < 128; i = i + 1) begin
        mem[i] <= 16'b0000000000000000;
      end
    end
  end

endmodule
